-- UndCC_Violation
library ieee;
use ieee.numeric_bit.all;
entity comp is
 port (a, b: in unsigned (7 downto 0);
 equal: out bit);
end comp;
architecture functional of comp is
begin
 process (a, b)
 begin
 if a = b then
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 equal <= '1';
 else
 equal <= '0';
 end if;
 end process;
end functional;
